module arm_verilog (OutD,OutC,A,D,Go,clk_in,reset_n);

input A,D,Go,clk_in,reset_n;
output OutD,OutC;
wire justWire;
reg justReg;

endmodule 
